LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX3_1 IS
PORT(
	ALU_B,RS_B,ADDR_B:IN STD_LOGIC;
	ALUOUT,RSOUT,ADDROUT:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	DBUS:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END MUX3_1;
ARCHITECTURE A OF MUX3_1 IS
BEGIN
	PROCESS
	BEGIN
		IF(ALU_B='0' AND RS_B='1' AND ADDR_B='1')THEN
			DBUS<=ALUOUT;
		ELSIF(ALU_B='1' AND RS_B='0' AND ADDR_B='1')THEN
			DBUS<=RSOUT;
		ELSIF(ALU_B='1' AND RS_B='1' AND ADDR_B='0')THEN
			DBUS<=ADDROUT;
		END IF;
	END PROCESS;
END A;
