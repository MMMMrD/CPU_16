LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ALU IS
PORT(
	X:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	Y:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	S2,S1,S0:IN STD_LOGIC;
	ALOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	ZF,CF:OUT STD_LOGIC
	);
END ALU;
ARCHITECTURE A OF ALU IS
SIGNAL XX,YY,TMP:STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
	PROCESS
	BEGIN
		IF(S2='0' AND S1='0' AND S0='0') THEN
			XX<='0'&X;
			YY<='0'&Y;
			TMP<=XX+YY;
			ALOUT<=TMP(7 DOWNTO 0);
			CF<=TMP(8);
			IF(TMP="100000000" OR TMP="000000000")THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S2='0' AND S1='0' AND S0='1') THEN
			XX<='0'&X;
			YY<='0'&Y;
			TMP<=XX-YY;
			ALOUT<=TMP(7 DOWNTO 0);
			CF<=TMP(8);
			IF(TMP="100000000" OR TMP="000000000")THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S2='0' AND S1='1' AND S0='0')THEN
			XX<='0'&X;
			TMP<=XX+1;
			ALOUT<=TMP(7 DOWNTO 0);
			CF<=TMP(8);
			IF(TMP="100000000" OR TMP="000000000")THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S2='0' AND S1='1' AND S0='1')THEN
			XX<='0'&X;
			TMP<=XX+1;
			ALOUT<=TMP(7 DOWNTO 0);
			CF<=TMP(8);
			IF(TMP="100000000" OR TMP="000000000")THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S2='1' AND S1='0' AND S0='0')THEN
			XX<='0'&X;
			YY<='0'&Y;
			TMP<=XX+YY;
			ALOUT<=TMP(7 DOWNTO 0);
			CF<=TMP(8);
			IF(TMP="100000000" OR TMP="000000000")THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S2='1' AND S1='0' AND S0='1')THEN
			XX<='0'&X;
			YY<='0'&Y;
			TMP<=XX+YY;
			ALOUT<=TMP(7 DOWNTO 0);
			CF<=TMP(8);
			IF(TMP="100000000" OR TMP="000000000")THEN
				ZF<='1';
			ELSE
				ZF<='0';
			END IF;
		ELSIF(S2='1' AND S1='1' AND S0='0')THEN
			ALOUT<=Y;
		END IF;
	END PROCESS;
END A;
			
			
	
