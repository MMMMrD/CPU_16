LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX4_2 IS
PORT(
	I9,I8:IN STD_LOGIC;
	X0,X1,X2,X3:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	W:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END MUX4_2;
ARCHITECTURE A OF MUX4_2 IS
BEGIN
	PROCESS
	BEGIN
		IF(I9='0' AND I8='0')THEN
			W<=X0;
		ELSIF(I9='0' AND I8='1')THEN
			W<=X1;
		ELSIF(I9='1' AND I8='0')THEN
			W<=X2;
		ELSE
			W<=X3;
		END IF;
	END PROCESS;
END A;
