LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX4_1 IS
PORT(
	I11,I10:IN STD_LOGIC;
	X0,X1,X2,X3:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	W:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END MUX4_1;
ARCHITECTURE A OF MUX4_1 IS
BEGIN
	PROCESS
	BEGIN
		IF(I11='0' AND I10='0')THEN
			W<=X0;
		ELSIF(I11='0' AND I10='1')THEN
			W<=X1;
		ELSIF(I11='1' AND I10='0')THEN
			W<=X2;
		ELSE
			W<=X3;
		END IF;
	END PROCESS;
END A;
