LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY ROM IS  
PORT( 
     DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0); 
     ADDR:IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
     CS:IN STD_LOGIC 
); 
END ROM; 
ARCHITECTURE A OF ROM IS 
BEGIN 
     DOUT<="1000000000000000" WHEN ADDR="00000000" AND CS='0' ELSE --0
           "1000000000000000" WHEN ADDR="00000001" AND CS='0' ELSE --1      
           "0000000000000000" WHEN ADDR="00000010" AND CS='0' ELSE --2        
           "1001001000000000" WHEN ADDR="00000011" AND CS='0' ELSE --3        
           "0000000000000000" WHEN ADDR="00000100" AND CS='0' ELSE --4         
           "1010000100000000" WHEN ADDR="00000101" AND CS='0' ELSE --5
           "1011000000000000" WHEN ADDR="00000110" AND CS='0' ELSE --6        
           "0000110100000000" WHEN ADDR="00000111" AND CS='0' ELSE --7        
           "1100011000000000" WHEN ADDR="00001000" AND CS='0' ELSE --8        
           "1101000100000000" WHEN ADDR="00001001" AND CS='0' ELSE --9        
           "1101000100000000" WHEN ADDR="00001010" AND CS='0' ELSE --10
           "1110000000000000" WHEN ADDR="00001011" AND CS='0' ELSE --11        
           "0000010100000000" WHEN ADDR="00001100" AND CS='0' ELSE --12        
           "1111100000000000" WHEN ADDR="00001101" AND CS='0' ELSE --13       
           "1110000000000000" WHEN ADDR="00001110" AND CS='0' ELSE --14       
           "0000110100000000" WHEN ADDR="00001111" AND CS='0' ELSE --15
           "0000110100000000" WHEN ADDR="00010000" AND CS='0' ELSE --16
           "0000110100000000" WHEN ADDR="00010001" AND CS='0' ELSE --17
           "0000110100000000" WHEN ADDR="00010010" AND CS='0' ELSE --18
           "0000110100000000" WHEN ADDR="00010011" AND CS='0' ELSE --19
           "0000110100000000" WHEN ADDR="00010100" AND CS='0' ELSE --20
           "0000110100000000" WHEN ADDR="00010101" AND CS='0' ELSE --21
           "0000110100000000" WHEN ADDR="00010110" AND CS='0' ELSE --22
           "0000110100000000" WHEN ADDR="00010111" AND CS='0' ELSE --23
           "0000110100000000" WHEN ADDR="00011000" AND CS='0' ELSE --24
           "0000110100000000" WHEN ADDR="00011001" AND CS='0' ELSE --25
           "0000110100000000" WHEN ADDR="00011010" AND CS='0' ELSE --26
           "0000110100000000" WHEN ADDR="00011011" AND CS='0' ELSE --27
           "0000110100000000" WHEN ADDR="00011100" AND CS='0' ELSE --28
           "0000110100000000" WHEN ADDR="00011101" AND CS='0' ELSE --29
           "0000110100000000" WHEN ADDR="00011110" AND CS='0' ELSE --30
           "0000110100000000" WHEN ADDR="00011111" AND CS='0' ELSE --31
           "0000110100000000" WHEN ADDR="00100000" AND CS='0' ELSE --32
           "1001000100000000" WHEN ADDR="00100001" AND CS='0' ELSE --33    
           "0000000100000000" WHEN ADDR="00100010" AND CS='0' ELSE --34       
           "1001001000000000" WHEN ADDR="00100011" AND CS='0' ELSE --35       
           "0000000000000000" WHEN ADDR="00100100" AND CS='0' ELSE --36        
           "1010000100000000" WHEN ADDR="00100101" AND CS='0' ELSE --37
           "1011000000000000" WHEN ADDR="00100110" AND CS='0' ELSE --38       
           "0000110100000000" WHEN ADDR="00100111" AND CS='0' ELSE --39       
           "1100011000000000" WHEN ADDR="00101000" AND CS='0' ELSE --40       
           "1101000100000000" WHEN ADDR="00101001" AND CS='0' ELSE --41       
           "1101000100000000" WHEN ADDR="00101010" AND CS='0' ELSE --42
           "1110000000000000" WHEN ADDR="00101011" AND CS='0' ELSE --43       
           "0000010100000000" WHEN ADDR="00101100" AND CS='0' ELSE --44       
           "1111100000000000" WHEN ADDR="00101101" AND CS='0' ELSE --45       
           "1110000000000000" WHEN ADDR="00101110" AND CS='0' ELSE --46
           "0000110100000000" WHEN ADDR="00101111" AND CS='0' ELSE --47
           "0000110100000000" WHEN ADDR="00110000" AND CS='0' ELSE --48
           "0000110100000000" WHEN ADDR="00110001" AND CS='0' ELSE --49
           "0000110100000000" WHEN ADDR="00110010" AND CS='0' ELSE --50
           "0000110100000000" WHEN ADDR="00110011" AND CS='0' ELSE --51
           "0000110100000000" WHEN ADDR="00110100" AND CS='0' ELSE --52
           "0000110100000000" WHEN ADDR="00110101" AND CS='0' ELSE --53
           "0000110100000000" WHEN ADDR="00110110" AND CS='0' ELSE --54
           "0000110100000000" WHEN ADDR="00110111" AND CS='0' ELSE --55
           "0000110100000000" WHEN ADDR="00111000" AND CS='0' ELSE --56
           "0000110100000000" WHEN ADDR="00111001" AND CS='0' ELSE --57
           "0000110100000000" WHEN ADDR="00111010" AND CS='0' ELSE --58
           "0000110100000000" WHEN ADDR="00111011" AND CS='0' ELSE --59
           "0000110100000000" WHEN ADDR="00111100" AND CS='0' ELSE --60
           "0000110100000000" WHEN ADDR="00111101" AND CS='0' ELSE --61
           "0000110100000000" WHEN ADDR="00111110" AND CS='0' ELSE --62
           "0000110100000000" WHEN ADDR="00111111" AND CS='0' ELSE --63
           "0000000000000000"; 
END A; 


