LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTROM IS 
PORT(
	ADDR:IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	UA:OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
	D:OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
);
END CONTROM;

ARCHITECTURE A OF CONTROM IS
SIGNAL DATAOUT:STD_LOGIC_VECTOR(25 DOWNTO 0);
BEGIN
	PROCESS(ADDR)
	BEGIN
		CASE ADDR IS
			WHEN "000000" => DATAOUT<="11010010001111110100000000";
			WHEN "000001" => DATAOUT<="11010010001111110100000000";
			WHEN "000010" => DATAOUT<="11010010001111110100000000";
			WHEN "000011" => DATAOUT<="11010010001111110100000000";
			WHEN "000100" => DATAOUT<="11010010001111110100000000";
			WHEN "000101" => DATAOUT<="11010010001111110100000000";
			WHEN "000110" => DATAOUT<="11010010001111110100000000";
			WHEN "000111" => DATAOUT<="11010010001111110100000000";
			WHEN "001000" => DATAOUT<="11010010001111110100000000";
			WHEN "001001" => DATAOUT<="11010010001111110100000000";
			WHEN "001010" => DATAOUT<="11010010001111110100000000";
			WHEN "001011" => DATAOUT<="11010010001111110100000000";
			WHEN "001100" => DATAOUT<="11010010001111110100000000";
			WHEN "001101" => DATAOUT<="11010010001111110100000000";
			WHEN "001110" => DATAOUT<="11010010001111110100000000";
			WHEN "001111" => DATAOUT<="11010010001111110100000000";
			WHEN "010000" => DATAOUT<="11010010001111110100000000";
			WHEN OTHERS => DATAOUT<="00000010001111111100000000";
		END CASE;
		UA(5 DOWNTO 0)<=DATAOUT(5 DOWNTO 0);
		D(19 DOWNTO 0)<=DATAOUT(23 DOWNTO 6);
	END PROCESS;
END A;
