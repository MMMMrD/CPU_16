LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MCOMMAND IS 
PORT(
	T2,T3,T4:IN STD_LOGIC;
	O:IN STD_LOGIC_VECTOR(19 DOWNTO 0);
	P1,P2:OUT STD_LOGIC;
	LOAD,LDPC,LDAR,LDIR,LDRI,RS_B,S2,S1,S0,ALU_B,RD_D,CS_D,RAM_B,CS_I,ADDR_B,SW_B,LED_B,LDPSW:OUT STD_LOGIC
);
END MCOMMAND;
ARCHITECTURE A OF MCOMMAND IS
SIGNAL DATAOUT:STD_LOGIC_VECTOR(19 DOWNTO 0);
BEGIN 
PROCESS(T2)
	BEGIN
		IF(T2'EVENT AND T2='1')THEN
			DATAOUT(19 DOWNTO 0)<=O(19 DOWNTO 0);
		END IF;
		P2<=O(0);
		P1<=O(1);
		LOAD<=O(19);
		LDPC<=O(18) AND T4;
		LDAR<=O(17) AND T3;
		LDIR<=O(16) AND T3;
		LDRI<=O(15) AND T4;
		RS_B<=O(13);
		S2<=O(12);
		S1<=O(11);
		S0<=O(10);
		ALU_B<=O(9);
		RD_D<=O(6);
		CS_D<=O(5);
		RAM_B<=O(4);
		CS_I<=O(3);
		ADDR_B<=O(2);
		SW_B<=O(8);
		LED_B<=O(7);
		LDPSW<=O(14) AND T4;
	END PROCESS;
END A;
